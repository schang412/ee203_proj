// Created by ihdl
module gen_stim (VDD, VSS, CLK_500K, VSTIM_P, VSTIM_N, MEASURE_PRESCALAR, DO_SAMPLE );
  input VDD;
  input VSS;
  input [3:0] MEASURE_PRESCALAR;
  input CLK_500K;
  output VSTIM_P, VSTIM_N, DO_SAMPLE;
  wire   N54, N55, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69,
         N70, N71, N72, N73, N74, N75, N76, n170, n250,
         rem_45_u_div_PartRem_30__2_, rem_45_u_div_PartRem_30__1_,
         rem_45_u_div_PartRem_29__3_, rem_45_u_div_PartRem_29__2_,
         rem_45_u_div_PartRem_29__1_, rem_45_u_div_PartRem_28__3_,
         rem_45_u_div_PartRem_28__2_, rem_45_u_div_PartRem_28__1_,
         rem_45_u_div_PartRem_27__3_, rem_45_u_div_PartRem_27__2_,
         rem_45_u_div_PartRem_27__1_, rem_45_u_div_PartRem_26__3_,
         rem_45_u_div_PartRem_26__2_, rem_45_u_div_PartRem_26__1_,
         rem_45_u_div_PartRem_25__3_, rem_45_u_div_PartRem_25__2_,
         rem_45_u_div_PartRem_25__1_, rem_45_u_div_PartRem_24__3_,
         rem_45_u_div_PartRem_24__2_, rem_45_u_div_PartRem_24__1_,
         rem_45_u_div_PartRem_23__3_, rem_45_u_div_PartRem_23__2_,
         rem_45_u_div_PartRem_23__1_, rem_45_u_div_PartRem_22__3_,
         rem_45_u_div_PartRem_22__2_, rem_45_u_div_PartRem_22__1_,
         rem_45_u_div_PartRem_21__3_, rem_45_u_div_PartRem_21__2_,
         rem_45_u_div_PartRem_21__1_, rem_45_u_div_PartRem_20__3_,
         rem_45_u_div_PartRem_20__2_, rem_45_u_div_PartRem_20__1_,
         rem_45_u_div_PartRem_19__3_, rem_45_u_div_PartRem_19__2_,
         rem_45_u_div_PartRem_19__1_, rem_45_u_div_PartRem_18__3_,
         rem_45_u_div_PartRem_18__2_, rem_45_u_div_PartRem_18__1_,
         rem_45_u_div_PartRem_17__3_, rem_45_u_div_PartRem_17__2_,
         rem_45_u_div_PartRem_17__1_, rem_45_u_div_PartRem_16__3_,
         rem_45_u_div_PartRem_16__2_, rem_45_u_div_PartRem_16__1_,
         rem_45_u_div_PartRem_15__3_, rem_45_u_div_PartRem_15__2_,
         rem_45_u_div_PartRem_15__1_, rem_45_u_div_PartRem_14__3_,
         rem_45_u_div_PartRem_14__2_, rem_45_u_div_PartRem_14__1_,
         rem_45_u_div_PartRem_13__3_, rem_45_u_div_PartRem_13__2_,
         rem_45_u_div_PartRem_13__1_, rem_45_u_div_PartRem_12__3_,
         rem_45_u_div_PartRem_12__2_, rem_45_u_div_PartRem_12__1_,
         rem_45_u_div_PartRem_11__3_, rem_45_u_div_PartRem_11__2_,
         rem_45_u_div_PartRem_11__1_, rem_45_u_div_PartRem_10__3_,
         rem_45_u_div_PartRem_10__2_, rem_45_u_div_PartRem_10__1_,
         rem_45_u_div_PartRem_9__3_, rem_45_u_div_PartRem_9__2_,
         rem_45_u_div_PartRem_9__1_, rem_45_u_div_PartRem_8__3_,
         rem_45_u_div_PartRem_8__2_, rem_45_u_div_PartRem_8__1_,
         rem_45_u_div_PartRem_7__3_, rem_45_u_div_PartRem_7__2_,
         rem_45_u_div_PartRem_7__1_, rem_45_u_div_PartRem_6__3_,
         rem_45_u_div_PartRem_6__2_, rem_45_u_div_PartRem_6__1_,
         rem_45_u_div_PartRem_5__3_, rem_45_u_div_PartRem_5__2_,
         rem_45_u_div_PartRem_5__1_, rem_45_u_div_PartRem_4__3_,
         rem_45_u_div_PartRem_4__2_, rem_45_u_div_PartRem_4__1_,
         rem_45_u_div_PartRem_3__3_, rem_45_u_div_PartRem_3__2_,
         rem_45_u_div_PartRem_3__1_, rem_45_u_div_PartRem_2__3_,
         rem_45_u_div_PartRem_2__2_, rem_45_u_div_PartRem_2__1_,
         rem_45_u_div_PartRem_1__3_, rem_45_u_div_PartRem_1__2_,
         rem_45_u_div_PartRem_1__1_, rem_45_u_div_CryTmp_30__2_,
         rem_45_u_div_CryTmp_30__1_, rem_45_u_div_CryTmp_29__3_,
         rem_45_u_div_CryTmp_29__2_, rem_45_u_div_CryTmp_29__1_,
         rem_45_u_div_CryTmp_28__4_, rem_45_u_div_CryTmp_28__3_,
         rem_45_u_div_CryTmp_28__2_, rem_45_u_div_CryTmp_28__1_,
         rem_45_u_div_CryTmp_27__4_, rem_45_u_div_CryTmp_27__3_,
         rem_45_u_div_CryTmp_27__2_, rem_45_u_div_CryTmp_27__1_,
         rem_45_u_div_CryTmp_26__4_, rem_45_u_div_CryTmp_26__3_,
         rem_45_u_div_CryTmp_26__2_, rem_45_u_div_CryTmp_26__1_,
         rem_45_u_div_CryTmp_25__4_, rem_45_u_div_CryTmp_25__3_,
         rem_45_u_div_CryTmp_25__2_, rem_45_u_div_CryTmp_25__1_,
         rem_45_u_div_CryTmp_24__4_, rem_45_u_div_CryTmp_24__3_,
         rem_45_u_div_CryTmp_24__2_, rem_45_u_div_CryTmp_24__1_,
         rem_45_u_div_CryTmp_23__4_, rem_45_u_div_CryTmp_23__3_,
         rem_45_u_div_CryTmp_23__2_, rem_45_u_div_CryTmp_23__1_,
         rem_45_u_div_CryTmp_22__4_, rem_45_u_div_CryTmp_22__3_,
         rem_45_u_div_CryTmp_22__2_, rem_45_u_div_CryTmp_22__1_,
         rem_45_u_div_CryTmp_21__4_, rem_45_u_div_CryTmp_21__3_,
         rem_45_u_div_CryTmp_21__2_, rem_45_u_div_CryTmp_21__1_,
         rem_45_u_div_CryTmp_20__4_, rem_45_u_div_CryTmp_20__3_,
         rem_45_u_div_CryTmp_20__2_, rem_45_u_div_CryTmp_20__1_,
         rem_45_u_div_CryTmp_19__4_, rem_45_u_div_CryTmp_19__3_,
         rem_45_u_div_CryTmp_19__2_, rem_45_u_div_CryTmp_19__1_,
         rem_45_u_div_CryTmp_18__4_, rem_45_u_div_CryTmp_18__3_,
         rem_45_u_div_CryTmp_18__2_, rem_45_u_div_CryTmp_18__1_,
         rem_45_u_div_CryTmp_17__4_, rem_45_u_div_CryTmp_17__3_,
         rem_45_u_div_CryTmp_17__2_, rem_45_u_div_CryTmp_17__1_,
         rem_45_u_div_CryTmp_16__4_, rem_45_u_div_CryTmp_16__3_,
         rem_45_u_div_CryTmp_16__2_, rem_45_u_div_CryTmp_16__1_,
         rem_45_u_div_CryTmp_15__4_, rem_45_u_div_CryTmp_15__3_,
         rem_45_u_div_CryTmp_15__2_, rem_45_u_div_CryTmp_15__1_,
         rem_45_u_div_CryTmp_14__4_, rem_45_u_div_CryTmp_14__3_,
         rem_45_u_div_CryTmp_14__2_, rem_45_u_div_CryTmp_14__1_,
         rem_45_u_div_CryTmp_13__4_, rem_45_u_div_CryTmp_13__3_,
         rem_45_u_div_CryTmp_13__2_, rem_45_u_div_CryTmp_13__1_,
         rem_45_u_div_CryTmp_12__4_, rem_45_u_div_CryTmp_12__3_,
         rem_45_u_div_CryTmp_12__2_, rem_45_u_div_CryTmp_12__1_,
         rem_45_u_div_CryTmp_11__4_, rem_45_u_div_CryTmp_11__3_,
         rem_45_u_div_CryTmp_11__2_, rem_45_u_div_CryTmp_11__1_,
         rem_45_u_div_CryTmp_10__4_, rem_45_u_div_CryTmp_10__3_,
         rem_45_u_div_CryTmp_10__2_, rem_45_u_div_CryTmp_10__1_,
         rem_45_u_div_CryTmp_9__4_, rem_45_u_div_CryTmp_9__3_,
         rem_45_u_div_CryTmp_9__2_, rem_45_u_div_CryTmp_9__1_,
         rem_45_u_div_CryTmp_8__4_, rem_45_u_div_CryTmp_8__3_,
         rem_45_u_div_CryTmp_8__2_, rem_45_u_div_CryTmp_8__1_,
         rem_45_u_div_CryTmp_7__4_, rem_45_u_div_CryTmp_7__3_,
         rem_45_u_div_CryTmp_7__2_, rem_45_u_div_CryTmp_7__1_,
         rem_45_u_div_CryTmp_6__4_, rem_45_u_div_CryTmp_6__3_,
         rem_45_u_div_CryTmp_6__2_, rem_45_u_div_CryTmp_6__1_,
         rem_45_u_div_CryTmp_5__4_, rem_45_u_div_CryTmp_5__3_,
         rem_45_u_div_CryTmp_5__2_, rem_45_u_div_CryTmp_5__1_,
         rem_45_u_div_CryTmp_4__4_, rem_45_u_div_CryTmp_4__3_,
         rem_45_u_div_CryTmp_4__2_, rem_45_u_div_CryTmp_4__1_,
         rem_45_u_div_CryTmp_3__4_, rem_45_u_div_CryTmp_3__3_,
         rem_45_u_div_CryTmp_3__2_, rem_45_u_div_CryTmp_3__1_,
         rem_45_u_div_CryTmp_2__4_, rem_45_u_div_CryTmp_2__3_,
         rem_45_u_div_CryTmp_2__2_, rem_45_u_div_CryTmp_2__1_,
         rem_45_u_div_CryTmp_1__4_, rem_45_u_div_CryTmp_1__3_,
         rem_45_u_div_CryTmp_1__2_, rem_45_u_div_CryTmp_1__1_,
         rem_45_u_div_CryTmp_0__4_, rem_45_u_div_CryTmp_0__3_,
         rem_45_u_div_CryTmp_0__2_, rem_45_u_div_SumTmp_30__1_,
         rem_45_u_div_SumTmp_29__2_, rem_45_u_div_SumTmp_29__1_,
         rem_45_u_div_SumTmp_28__3_, rem_45_u_div_SumTmp_28__2_,
         rem_45_u_div_SumTmp_28__1_, rem_45_u_div_SumTmp_27__3_,
         rem_45_u_div_SumTmp_27__2_, rem_45_u_div_SumTmp_27__1_,
         rem_45_u_div_SumTmp_26__3_, rem_45_u_div_SumTmp_26__2_,
         rem_45_u_div_SumTmp_26__1_, rem_45_u_div_SumTmp_25__3_,
         rem_45_u_div_SumTmp_25__2_, rem_45_u_div_SumTmp_25__1_,
         rem_45_u_div_SumTmp_24__3_, rem_45_u_div_SumTmp_24__2_,
         rem_45_u_div_SumTmp_24__1_, rem_45_u_div_SumTmp_23__3_,
         rem_45_u_div_SumTmp_23__2_, rem_45_u_div_SumTmp_23__1_,
         rem_45_u_div_SumTmp_22__3_, rem_45_u_div_SumTmp_22__2_,
         rem_45_u_div_SumTmp_22__1_, rem_45_u_div_SumTmp_21__3_,
         rem_45_u_div_SumTmp_21__2_, rem_45_u_div_SumTmp_21__1_,
         rem_45_u_div_SumTmp_20__3_, rem_45_u_div_SumTmp_20__2_,
         rem_45_u_div_SumTmp_20__1_, rem_45_u_div_SumTmp_19__3_,
         rem_45_u_div_SumTmp_19__2_, rem_45_u_div_SumTmp_19__1_,
         rem_45_u_div_SumTmp_18__3_, rem_45_u_div_SumTmp_18__2_,
         rem_45_u_div_SumTmp_18__1_, rem_45_u_div_SumTmp_17__3_,
         rem_45_u_div_SumTmp_17__2_, rem_45_u_div_SumTmp_17__1_,
         rem_45_u_div_SumTmp_16__3_, rem_45_u_div_SumTmp_16__2_,
         rem_45_u_div_SumTmp_16__1_, rem_45_u_div_SumTmp_15__3_,
         rem_45_u_div_SumTmp_15__2_, rem_45_u_div_SumTmp_15__1_,
         rem_45_u_div_SumTmp_14__3_, rem_45_u_div_SumTmp_14__2_,
         rem_45_u_div_SumTmp_14__1_, rem_45_u_div_SumTmp_13__3_,
         rem_45_u_div_SumTmp_13__2_, rem_45_u_div_SumTmp_13__1_,
         rem_45_u_div_SumTmp_12__3_, rem_45_u_div_SumTmp_12__2_,
         rem_45_u_div_SumTmp_12__1_, rem_45_u_div_SumTmp_11__3_,
         rem_45_u_div_SumTmp_11__2_, rem_45_u_div_SumTmp_11__1_,
         rem_45_u_div_SumTmp_10__3_, rem_45_u_div_SumTmp_10__2_,
         rem_45_u_div_SumTmp_10__1_, rem_45_u_div_SumTmp_9__3_,
         rem_45_u_div_SumTmp_9__2_, rem_45_u_div_SumTmp_9__1_,
         rem_45_u_div_SumTmp_8__3_, rem_45_u_div_SumTmp_8__2_,
         rem_45_u_div_SumTmp_8__1_, rem_45_u_div_SumTmp_7__3_,
         rem_45_u_div_SumTmp_7__2_, rem_45_u_div_SumTmp_7__1_,
         rem_45_u_div_SumTmp_6__3_, rem_45_u_div_SumTmp_6__2_,
         rem_45_u_div_SumTmp_6__1_, rem_45_u_div_SumTmp_5__3_,
         rem_45_u_div_SumTmp_5__2_, rem_45_u_div_SumTmp_5__1_,
         rem_45_u_div_SumTmp_4__3_, rem_45_u_div_SumTmp_4__2_,
         rem_45_u_div_SumTmp_4__1_, rem_45_u_div_SumTmp_3__3_,
         rem_45_u_div_SumTmp_3__2_, rem_45_u_div_SumTmp_3__1_,
         rem_45_u_div_SumTmp_2__3_, rem_45_u_div_SumTmp_2__2_,
         rem_45_u_div_SumTmp_2__1_, rem_45_u_div_SumTmp_1__3_,
         rem_45_u_div_SumTmp_1__2_, rem_45_u_div_SumTmp_1__1_,
         rem_45_u_div_SumTmp_0__3_, rem_45_u_div_SumTmp_0__2_,
         rem_45_u_div_SumTmp_0__1_, n43, n440, n47, n48, n49, n50, n51, n52,
         n53, n540, n550, n56, n57, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n229, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n247, n248, n249, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n320, n321, n323, n325, n326, n327, n328, n330,
         n331, n333, n335, n336, n337, n338, n341, n342, n344, n346, n347,
         n348, n350, n351, n353, n354, n356, n357, n359, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n413, n414,
         n415, n416, n417, n418, n420, n421, n422, n423, n424, n425, n426,
         n432, n433, n434, n436, n437, n438, n439, n441;

  AO22_F U61 ( .A1(rem_45_u_div_SumTmp_1__1_), .A2(n191), .B1(n257), .B2(
        rem_45_u_div_PartRem_2__1_), .Z(rem_45_u_div_PartRem_1__2_) );
  AO22_F U65 ( .A1(rem_45_u_div_SumTmp_1__2_), .A2(n191), .B1(n257), .B2(
        rem_45_u_div_PartRem_2__2_), .Z(rem_45_u_div_PartRem_1__3_) );
  AO22_F U66 ( .A1(rem_45_u_div_SumTmp_2__1_), .A2(n192), .B1(n259), .B2(
        rem_45_u_div_PartRem_3__1_), .Z(rem_45_u_div_PartRem_2__2_) );
  AO22_F U75 ( .A1(rem_45_u_div_SumTmp_2__2_), .A2(n192), .B1(n259), .B2(
        rem_45_u_div_PartRem_3__2_), .Z(rem_45_u_div_PartRem_2__3_) );
  AO22_F U76 ( .A1(rem_45_u_div_SumTmp_3__1_), .A2(n264), .B1(n193), .B2(
        rem_45_u_div_PartRem_4__1_), .Z(rem_45_u_div_PartRem_3__2_) );
  AO21_I U78 ( .A1(n194), .A2(n438), .B(n48), .Z(n266) );
  AO21_I U81 ( .A1(n259), .A2(rem_45_u_div_PartRem_3__3_), .B(
        rem_45_u_div_CryTmp_1__4_), .Z(n267) );
  AO22_F U82 ( .A1(rem_45_u_div_SumTmp_3__2_), .A2(n264), .B1(n193), .B2(
        rem_45_u_div_PartRem_4__2_), .Z(rem_45_u_div_PartRem_3__3_) );
  AO22_F U83 ( .A1(rem_45_u_div_SumTmp_4__1_), .A2(n194), .B1(n265), .B2(
        rem_45_u_div_PartRem_5__1_), .Z(rem_45_u_div_PartRem_4__2_) );
  AO21_I U88 ( .A1(n193), .A2(rem_45_u_div_PartRem_4__3_), .B(
        rem_45_u_div_CryTmp_2__4_), .Z(n271) );
  AO22_F U89 ( .A1(rem_45_u_div_SumTmp_4__2_), .A2(n194), .B1(n265), .B2(
        rem_45_u_div_PartRem_5__2_), .Z(rem_45_u_div_PartRem_4__3_) );
  AO22_F U90 ( .A1(rem_45_u_div_SumTmp_5__1_), .A2(n195), .B1(n268), .B2(
        rem_45_u_div_PartRem_6__1_), .Z(rem_45_u_div_PartRem_5__2_) );
  AO21_I U92 ( .A1(n273), .A2(n438), .B(n50), .Z(n272) );
  AO22_F U97 ( .A1(rem_45_u_div_SumTmp_5__2_), .A2(n195), .B1(n268), .B2(
        rem_45_u_div_PartRem_6__2_), .Z(rem_45_u_div_PartRem_5__3_) );
  AO22_F U98 ( .A1(rem_45_u_div_SumTmp_6__1_), .A2(n273), .B1(n196), .B2(
        rem_45_u_div_PartRem_7__1_), .Z(rem_45_u_div_PartRem_6__2_) );
  AO21_I U103 ( .A1(n268), .A2(rem_45_u_div_PartRem_6__3_), .B(
        rem_45_u_div_CryTmp_4__4_), .Z(n278) );
  AO22_F U104 ( .A1(rem_45_u_div_SumTmp_6__2_), .A2(n273), .B1(n196), .B2(
        rem_45_u_div_PartRem_7__2_), .Z(rem_45_u_div_PartRem_6__3_) );
  AO22_F U105 ( .A1(rem_45_u_div_SumTmp_7__1_), .A2(n197), .B1(n276), .B2(
        rem_45_u_div_PartRem_8__1_), .Z(rem_45_u_div_PartRem_7__2_) );
  AO21_I U107 ( .A1(n207), .A2(n438), .B(n52), .Z(n280) );
  AO21_I U110 ( .A1(n196), .A2(rem_45_u_div_PartRem_7__3_), .B(
        rem_45_u_div_CryTmp_5__4_), .Z(n281) );
  AO22_F U111 ( .A1(rem_45_u_div_SumTmp_7__2_), .A2(n197), .B1(n276), .B2(
        rem_45_u_div_PartRem_8__2_), .Z(rem_45_u_div_PartRem_7__3_) );
  AO22_F U112 ( .A1(rem_45_u_div_SumTmp_8__1_), .A2(n207), .B1(n279), .B2(
        rem_45_u_div_PartRem_9__1_), .Z(rem_45_u_div_PartRem_8__2_) );
  AO22_F U119 ( .A1(rem_45_u_div_SumTmp_8__2_), .A2(n207), .B1(n279), .B2(
        rem_45_u_div_PartRem_9__2_), .Z(rem_45_u_div_PartRem_8__3_) );
  AO22_F U120 ( .A1(rem_45_u_div_SumTmp_9__1_), .A2(n285), .B1(n208), .B2(
        rem_45_u_div_PartRem_10__1_), .Z(rem_45_u_div_PartRem_9__2_) );
  AO21_I U125 ( .A1(n279), .A2(rem_45_u_div_PartRem_9__3_), .B(
        rem_45_u_div_CryTmp_7__4_), .Z(n288) );
  AO22_F U126 ( .A1(rem_45_u_div_SumTmp_9__2_), .A2(n285), .B1(n208), .B2(
        rem_45_u_div_PartRem_10__2_), .Z(rem_45_u_div_PartRem_9__3_) );
  AO22_F U127 ( .A1(rem_45_u_div_SumTmp_10__1_), .A2(n210), .B1(n286), .B2(
        rem_45_u_div_PartRem_11__1_), .Z(rem_45_u_div_PartRem_10__2_) );
  AO21_I U132 ( .A1(n208), .A2(rem_45_u_div_PartRem_10__3_), .B(
        rem_45_u_div_CryTmp_8__4_), .Z(n292) );
  AO22_F U133 ( .A1(rem_45_u_div_SumTmp_10__2_), .A2(n210), .B1(n286), .B2(
        rem_45_u_div_PartRem_11__2_), .Z(rem_45_u_div_PartRem_10__3_) );
  AO22_F U134 ( .A1(rem_45_u_div_SumTmp_11__1_), .A2(n212), .B1(n289), .B2(
        rem_45_u_div_PartRem_12__1_), .Z(rem_45_u_div_PartRem_11__2_) );
  AO21_I U136 ( .A1(n294), .A2(n438), .B(n550), .Z(n293) );
  AO22_F U141 ( .A1(rem_45_u_div_SumTmp_11__2_), .A2(n212), .B1(n289), .B2(
        rem_45_u_div_PartRem_12__2_), .Z(rem_45_u_div_PartRem_11__3_) );
  AO22_F U142 ( .A1(rem_45_u_div_SumTmp_12__1_), .A2(n294), .B1(n214), .B2(
        rem_45_u_div_PartRem_13__1_), .Z(rem_45_u_div_PartRem_12__2_) );
  AO21_I U147 ( .A1(n289), .A2(rem_45_u_div_PartRem_12__3_), .B(
        rem_45_u_div_CryTmp_10__4_), .Z(n299) );
  AO22_F U148 ( .A1(rem_45_u_div_SumTmp_12__2_), .A2(n294), .B1(n214), .B2(
        rem_45_u_div_PartRem_13__2_), .Z(rem_45_u_div_PartRem_12__3_) );
  AO22_F U149 ( .A1(rem_45_u_div_SumTmp_13__1_), .A2(n215), .B1(n297), .B2(
        rem_45_u_div_PartRem_14__1_), .Z(rem_45_u_div_PartRem_13__2_) );
  AO21_I U154 ( .A1(n214), .A2(rem_45_u_div_PartRem_13__3_), .B(
        rem_45_u_div_CryTmp_11__4_), .Z(n303) );
  AO22_F U155 ( .A1(rem_45_u_div_SumTmp_13__2_), .A2(n215), .B1(n297), .B2(
        rem_45_u_div_PartRem_14__2_), .Z(rem_45_u_div_PartRem_13__3_) );
  AO22_F U156 ( .A1(rem_45_u_div_SumTmp_14__1_), .A2(n217), .B1(n301), .B2(
        rem_45_u_div_PartRem_15__1_), .Z(rem_45_u_div_PartRem_14__2_) );
  AO22_F U163 ( .A1(rem_45_u_div_SumTmp_14__2_), .A2(n217), .B1(n301), .B2(
        rem_45_u_div_PartRem_15__2_), .Z(rem_45_u_div_PartRem_14__3_) );
  AO22_F U164 ( .A1(rem_45_u_div_SumTmp_15__1_), .A2(n307), .B1(n219), .B2(
        rem_45_u_div_PartRem_16__1_), .Z(rem_45_u_div_PartRem_15__2_) );
  AO21_I U169 ( .A1(n301), .A2(rem_45_u_div_PartRem_15__3_), .B(
        rem_45_u_div_CryTmp_13__4_), .Z(n310) );
  AO22_F U170 ( .A1(rem_45_u_div_SumTmp_15__2_), .A2(n307), .B1(n219), .B2(
        rem_45_u_div_PartRem_16__2_), .Z(rem_45_u_div_PartRem_15__3_) );
  AO22_F U171 ( .A1(rem_45_u_div_SumTmp_16__1_), .A2(n221), .B1(n308), .B2(
        rem_45_u_div_PartRem_17__1_), .Z(rem_45_u_div_PartRem_16__2_) );
  AO21_I U176 ( .A1(n219), .A2(rem_45_u_div_PartRem_16__3_), .B(
        rem_45_u_div_CryTmp_14__4_), .Z(n313) );
  AO22_F U177 ( .A1(rem_45_u_div_SumTmp_16__2_), .A2(n221), .B1(n308), .B2(
        rem_45_u_div_PartRem_17__2_), .Z(rem_45_u_div_PartRem_16__3_) );
  AO22_F U178 ( .A1(rem_45_u_div_SumTmp_17__1_), .A2(n223), .B1(n311), .B2(
        rem_45_u_div_PartRem_18__1_), .Z(rem_45_u_div_PartRem_17__2_) );
  AO22_F U185 ( .A1(rem_45_u_div_SumTmp_17__2_), .A2(n223), .B1(n311), .B2(
        rem_45_u_div_PartRem_18__2_), .Z(rem_45_u_div_PartRem_17__3_) );
  AO22_F U186 ( .A1(rem_45_u_div_SumTmp_18__1_), .A2(n317), .B1(n225), .B2(
        rem_45_u_div_PartRem_19__1_), .Z(rem_45_u_div_PartRem_18__2_) );
  AO21_I U191 ( .A1(n311), .A2(rem_45_u_div_PartRem_18__3_), .B(
        rem_45_u_div_CryTmp_16__4_), .Z(n320) );
  AO22_F U192 ( .A1(rem_45_u_div_SumTmp_18__2_), .A2(n317), .B1(n225), .B2(
        rem_45_u_div_PartRem_19__2_), .Z(rem_45_u_div_PartRem_18__3_) );
  AO22_F U193 ( .A1(rem_45_u_div_SumTmp_19__1_), .A2(n227), .B1(n318), .B2(
        rem_45_u_div_PartRem_20__1_), .Z(rem_45_u_div_PartRem_19__2_) );
  AO21_I U198 ( .A1(n225), .A2(rem_45_u_div_PartRem_19__3_), .B(
        rem_45_u_div_CryTmp_17__4_), .Z(n323) );
  AO22_F U199 ( .A1(rem_45_u_div_SumTmp_19__2_), .A2(n227), .B1(n318), .B2(
        rem_45_u_div_PartRem_20__2_), .Z(rem_45_u_div_PartRem_19__3_) );
  AO22_F U200 ( .A1(rem_45_u_div_SumTmp_20__1_), .A2(n229), .B1(n321), .B2(
        rem_45_u_div_PartRem_21__1_), .Z(rem_45_u_div_PartRem_20__2_) );
  AO22_F U207 ( .A1(rem_45_u_div_SumTmp_20__2_), .A2(n229), .B1(n321), .B2(
        rem_45_u_div_PartRem_21__2_), .Z(rem_45_u_div_PartRem_20__3_) );
  AO22_F U208 ( .A1(rem_45_u_div_SumTmp_21__1_), .A2(n325), .B1(n231), .B2(
        rem_45_u_div_PartRem_22__1_), .Z(rem_45_u_div_PartRem_21__2_) );
  AO21_I U213 ( .A1(n321), .A2(rem_45_u_div_PartRem_21__3_), .B(
        rem_45_u_div_CryTmp_19__4_), .Z(n330) );
  AO22_F U214 ( .A1(rem_45_u_div_SumTmp_21__2_), .A2(n325), .B1(n231), .B2(
        rem_45_u_div_PartRem_22__2_), .Z(rem_45_u_div_PartRem_21__3_) );
  AO22_F U215 ( .A1(rem_45_u_div_SumTmp_22__1_), .A2(n232), .B1(n328), .B2(
        rem_45_u_div_PartRem_23__1_), .Z(rem_45_u_div_PartRem_22__2_) );
  AO21_I U220 ( .A1(n231), .A2(rem_45_u_div_PartRem_22__3_), .B(
        rem_45_u_div_CryTmp_20__4_), .Z(n333) );
  AO22_F U221 ( .A1(rem_45_u_div_SumTmp_22__2_), .A2(n232), .B1(n328), .B2(
        rem_45_u_div_PartRem_23__2_), .Z(rem_45_u_div_PartRem_22__3_) );
  AO22_F U222 ( .A1(rem_45_u_div_SumTmp_23__1_), .A2(n233), .B1(n331), .B2(
        rem_45_u_div_PartRem_24__1_), .Z(rem_45_u_div_PartRem_23__2_) );
  AO22_F U229 ( .A1(rem_45_u_div_SumTmp_23__2_), .A2(n233), .B1(n331), .B2(
        rem_45_u_div_PartRem_24__2_), .Z(rem_45_u_div_PartRem_23__3_) );
  AO22_F U230 ( .A1(rem_45_u_div_SumTmp_24__1_), .A2(n335), .B1(n234), .B2(
        rem_45_u_div_PartRem_25__1_), .Z(rem_45_u_div_PartRem_24__2_) );
  AO21_I U235 ( .A1(n331), .A2(rem_45_u_div_PartRem_24__3_), .B(
        rem_45_u_div_CryTmp_22__4_), .Z(n341) );
  AO22_F U236 ( .A1(rem_45_u_div_SumTmp_24__2_), .A2(n335), .B1(n234), .B2(
        rem_45_u_div_PartRem_25__2_), .Z(rem_45_u_div_PartRem_24__3_) );
  AO22_F U237 ( .A1(rem_45_u_div_SumTmp_25__1_), .A2(n235), .B1(n338), .B2(
        rem_45_u_div_PartRem_26__1_), .Z(rem_45_u_div_PartRem_25__2_) );
  AO21_I U242 ( .A1(n234), .A2(rem_45_u_div_PartRem_25__3_), .B(
        rem_45_u_div_CryTmp_23__4_), .Z(n344) );
  AO22_F U243 ( .A1(rem_45_u_div_SumTmp_25__2_), .A2(n235), .B1(n338), .B2(
        rem_45_u_div_PartRem_26__2_), .Z(rem_45_u_div_PartRem_25__3_) );
  AO22_F U244 ( .A1(rem_45_u_div_SumTmp_26__1_), .A2(n236), .B1(n342), .B2(
        rem_45_u_div_PartRem_27__1_), .Z(rem_45_u_div_PartRem_26__2_) );
  AO22_F U251 ( .A1(rem_45_u_div_SumTmp_26__2_), .A2(n236), .B1(n342), .B2(
        rem_45_u_div_PartRem_27__2_), .Z(rem_45_u_div_PartRem_26__3_) );
  AO22_F U252 ( .A1(rem_45_u_div_SumTmp_27__1_), .A2(n346), .B1(n237), .B2(
        rem_45_u_div_PartRem_28__1_), .Z(rem_45_u_div_PartRem_27__2_) );
  AO21_I U257 ( .A1(n342), .A2(rem_45_u_div_PartRem_27__3_), .B(
        rem_45_u_div_CryTmp_25__4_), .Z(n350) );
  AO22_F U258 ( .A1(rem_45_u_div_SumTmp_27__2_), .A2(n346), .B1(n237), .B2(
        rem_45_u_div_PartRem_28__2_), .Z(rem_45_u_div_PartRem_27__3_) );
  AO22_F U259 ( .A1(rem_45_u_div_SumTmp_28__1_), .A2(
        rem_45_u_div_CryTmp_28__4_), .B1(rem_45_u_div_PartRem_29__1_), .B2(
        n238), .Z(rem_45_u_div_PartRem_28__2_) );
  AO21_I U264 ( .A1(n237), .A2(rem_45_u_div_PartRem_28__3_), .B(
        rem_45_u_div_CryTmp_26__4_), .Z(n353) );
  AO22_F U265 ( .A1(rem_45_u_div_SumTmp_28__2_), .A2(
        rem_45_u_div_CryTmp_28__4_), .B1(rem_45_u_div_PartRem_29__2_), .B2(
        n238), .Z(rem_45_u_div_PartRem_28__3_) );
  AO22_F U266 ( .A1(rem_45_u_div_SumTmp_29__1_), .A2(n239), .B1(
        rem_45_u_div_PartRem_30__1_), .B2(n351), .Z(
        rem_45_u_div_PartRem_29__2_) );
  AO22_F U273 ( .A1(rem_45_u_div_SumTmp_29__2_), .A2(n239), .B1(
        rem_45_u_div_PartRem_30__2_), .B2(n351), .Z(
        rem_45_u_div_PartRem_29__3_) );
  XNOR2_C U283 ( .A(n224), .B(n362), .Z(n363) );
  XNOR2_C U286 ( .A(n364), .B(n57), .Z(n365) );
  XNOR2_C U289 ( .A(n220), .B(n366), .Z(n367) );
  XNOR2_C U292 ( .A(n368), .B(n424), .Z(n369) );
  XNOR2_C U295 ( .A(n216), .B(n370), .Z(n371) );
  XNOR2_C U298 ( .A(n372), .B(n550), .Z(n373) );
  XNOR2_C U301 ( .A(n213), .B(n374), .Z(n375) );
  XNOR2_C U304 ( .A(n376), .B(n423), .Z(n377) );
  XNOR2_C U307 ( .A(n209), .B(n378), .Z(n379) );
  XNOR2_C U310 ( .A(n381), .B(n52), .Z(n382) );
  XNOR2_C U313 ( .A(n198), .B(n383), .Z(n384) );
  XNOR2_C U316 ( .A(n385), .B(n50), .Z(n386) );
  XNOR2_C U319 ( .A(n206), .B(n387), .Z(n388) );
  XNOR2_C U322 ( .A(n389), .B(n48), .Z(n390) );
  XNOR2_C U325 ( .A(n201), .B(n391), .Z(n392) );
  XNOR2_C U331 ( .A(n204), .B(n205), .Z(n395) );
  AO21_I U345 ( .A1(n413), .A2(n211), .B(n414), .Z(n251) );
  INVERTBAL_H U363 ( .A(n256), .Z(n190) );
  INVERTBAL_H U364 ( .A(n257), .Z(n191) );
  INVERTBAL_H U365 ( .A(n259), .Z(n192) );
  INVERTBAL_H U366 ( .A(n264), .Z(n193) );
  INVERTBAL_H U367 ( .A(n265), .Z(n194) );
  INVERTBAL_H U368 ( .A(n268), .Z(n195) );
  INVERTBAL_H U369 ( .A(n273), .Z(n196) );
  INVERTBAL_H U370 ( .A(n276), .Z(n197) );
  INVERTBAL_H U372 ( .A(n436), .Z(n199) );
  INVERTBAL_H U373 ( .A(n408), .Z(n200) );
  INVERTBAL_H U376 ( .A(n247), .Z(n203) );
  INVERTBAL_H U380 ( .A(n279), .Z(n207) );
  INVERTBAL_H U381 ( .A(n285), .Z(n208) );
  INVERTBAL_H U383 ( .A(n286), .Z(n210) );
  INVERTBAL_H U385 ( .A(n289), .Z(n212) );
  INVERTBAL_H U387 ( .A(n294), .Z(n214) );
  INVERTBAL_H U388 ( .A(n297), .Z(n215) );
  INVERTBAL_H U390 ( .A(n301), .Z(n217) );
  INVERTBAL_H U392 ( .A(n307), .Z(n219) );
  INVERTBAL_H U394 ( .A(n308), .Z(n221) );
  INVERTBAL_H U396 ( .A(n311), .Z(n223) );
  INVERTBAL_H U398 ( .A(n317), .Z(n225) );
  INVERTBAL_H U400 ( .A(n318), .Z(n227) );
  INVERTBAL_H U402 ( .A(n321), .Z(n229) );
  INVERTBAL_H U404 ( .A(n325), .Z(n231) );
  INVERTBAL_H U405 ( .A(n328), .Z(n232) );
  INVERTBAL_H U406 ( .A(n331), .Z(n233) );
  INVERTBAL_H U407 ( .A(n335), .Z(n234) );
  INVERTBAL_H U408 ( .A(n338), .Z(n235) );
  INVERTBAL_H U409 ( .A(n342), .Z(n236) );
  INVERTBAL_H U410 ( .A(n346), .Z(n237) );
  INVERTBAL_H U411 ( .A(rem_45_u_div_CryTmp_28__4_), .Z(n238) );
  INVERTBAL_H U412 ( .A(n351), .Z(n239) );
  INVERTBAL_H U413 ( .A(n354), .Z(n240) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_0_1 ( .A(rem_45_u_div_PartRem_1__1_), .B(
        n243), .CIN(n203), .COUT(rem_45_u_div_CryTmp_0__2_), .SUM(
        rem_45_u_div_SumTmp_0__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_5_1 ( .A(rem_45_u_div_PartRem_6__1_), .B(
        n243), .CIN(rem_45_u_div_CryTmp_5__1_), .COUT(
        rem_45_u_div_CryTmp_5__2_), .SUM(rem_45_u_div_SumTmp_5__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_0_2 ( .A(rem_45_u_div_PartRem_1__2_), .B(
        n242), .CIN(rem_45_u_div_CryTmp_0__2_), .COUT(
        rem_45_u_div_CryTmp_0__3_), .SUM(rem_45_u_div_SumTmp_0__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_7_1 ( .A(rem_45_u_div_PartRem_8__1_), .B(
        n243), .CIN(rem_45_u_div_CryTmp_7__1_), .COUT(
        rem_45_u_div_CryTmp_7__2_), .SUM(rem_45_u_div_SumTmp_7__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_8_1 ( .A(rem_45_u_div_PartRem_9__1_), .B(
        n243), .CIN(rem_45_u_div_CryTmp_8__1_), .COUT(
        rem_45_u_div_CryTmp_8__2_), .SUM(rem_45_u_div_SumTmp_8__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_1_2 ( .A(rem_45_u_div_PartRem_2__2_), .B(
        n242), .CIN(rem_45_u_div_CryTmp_1__2_), .COUT(
        rem_45_u_div_CryTmp_1__3_), .SUM(rem_45_u_div_SumTmp_1__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_1_1 ( .A(rem_45_u_div_PartRem_2__1_), .B(
        n243), .CIN(rem_45_u_div_CryTmp_1__1_), .COUT(
        rem_45_u_div_CryTmp_1__2_), .SUM(rem_45_u_div_SumTmp_1__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_2_2 ( .A(rem_45_u_div_PartRem_3__2_), .B(
        n242), .CIN(rem_45_u_div_CryTmp_2__2_), .COUT(
        rem_45_u_div_CryTmp_2__3_), .SUM(rem_45_u_div_SumTmp_2__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_2_1 ( .A(rem_45_u_div_PartRem_3__1_), .B(
        n243), .CIN(rem_45_u_div_CryTmp_2__1_), .COUT(
        rem_45_u_div_CryTmp_2__2_), .SUM(rem_45_u_div_SumTmp_2__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_3_2 ( .A(rem_45_u_div_PartRem_4__2_), .B(
        n242), .CIN(rem_45_u_div_CryTmp_3__2_), .COUT(
        rem_45_u_div_CryTmp_3__3_), .SUM(rem_45_u_div_SumTmp_3__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_3_1 ( .A(rem_45_u_div_PartRem_4__1_), .B(
        n243), .CIN(rem_45_u_div_CryTmp_3__1_), .COUT(
        rem_45_u_div_CryTmp_3__2_), .SUM(rem_45_u_div_SumTmp_3__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_4_2 ( .A(rem_45_u_div_PartRem_5__2_), .B(
        n242), .CIN(rem_45_u_div_CryTmp_4__2_), .COUT(
        rem_45_u_div_CryTmp_4__3_), .SUM(rem_45_u_div_SumTmp_4__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_4_1 ( .A(rem_45_u_div_PartRem_5__1_), .B(
        n243), .CIN(rem_45_u_div_CryTmp_4__1_), .COUT(
        rem_45_u_div_CryTmp_4__2_), .SUM(rem_45_u_div_SumTmp_4__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_5_2 ( .A(rem_45_u_div_PartRem_6__2_), .B(
        n242), .CIN(rem_45_u_div_CryTmp_5__2_), .COUT(
        rem_45_u_div_CryTmp_5__3_), .SUM(rem_45_u_div_SumTmp_5__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_6_2 ( .A(rem_45_u_div_PartRem_7__2_), .B(
        n242), .CIN(rem_45_u_div_CryTmp_6__2_), .COUT(
        rem_45_u_div_CryTmp_6__3_), .SUM(rem_45_u_div_SumTmp_6__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_6_1 ( .A(rem_45_u_div_PartRem_7__1_), .B(
        n243), .CIN(rem_45_u_div_CryTmp_6__1_), .COUT(
        rem_45_u_div_CryTmp_6__2_), .SUM(rem_45_u_div_SumTmp_6__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_7_2 ( .A(rem_45_u_div_PartRem_8__2_), .B(
        n242), .CIN(rem_45_u_div_CryTmp_7__2_), .COUT(
        rem_45_u_div_CryTmp_7__3_), .SUM(rem_45_u_div_SumTmp_7__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_8_2 ( .A(rem_45_u_div_PartRem_9__2_), .B(
        n242), .CIN(rem_45_u_div_CryTmp_8__2_), .COUT(
        rem_45_u_div_CryTmp_8__3_), .SUM(rem_45_u_div_SumTmp_8__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_9_2 ( .A(rem_45_u_div_PartRem_10__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_9__2_), .COUT(
        rem_45_u_div_CryTmp_9__3_), .SUM(rem_45_u_div_SumTmp_9__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_9_1 ( .A(rem_45_u_div_PartRem_10__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_9__1_), .COUT(
        rem_45_u_div_CryTmp_9__2_), .SUM(rem_45_u_div_SumTmp_9__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_10_2 ( .A(rem_45_u_div_PartRem_11__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_10__2_), .COUT(
        rem_45_u_div_CryTmp_10__3_), .SUM(rem_45_u_div_SumTmp_10__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_10_1 ( .A(rem_45_u_div_PartRem_11__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_10__1_), .COUT(
        rem_45_u_div_CryTmp_10__2_), .SUM(rem_45_u_div_SumTmp_10__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_11_2 ( .A(rem_45_u_div_PartRem_12__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_11__2_), .COUT(
        rem_45_u_div_CryTmp_11__3_), .SUM(rem_45_u_div_SumTmp_11__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_11_1 ( .A(rem_45_u_div_PartRem_12__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_11__1_), .COUT(
        rem_45_u_div_CryTmp_11__2_), .SUM(rem_45_u_div_SumTmp_11__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_12_2 ( .A(rem_45_u_div_PartRem_13__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_12__2_), .COUT(
        rem_45_u_div_CryTmp_12__3_), .SUM(rem_45_u_div_SumTmp_12__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_12_1 ( .A(rem_45_u_div_PartRem_13__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_12__1_), .COUT(
        rem_45_u_div_CryTmp_12__2_), .SUM(rem_45_u_div_SumTmp_12__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_25_2 ( .A(rem_45_u_div_PartRem_26__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_25__2_), .COUT(
        rem_45_u_div_CryTmp_25__3_), .SUM(rem_45_u_div_SumTmp_25__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_25_1 ( .A(rem_45_u_div_PartRem_26__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_25__1_), .COUT(
        rem_45_u_div_CryTmp_25__2_), .SUM(rem_45_u_div_SumTmp_25__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_4_3 ( .A(rem_45_u_div_PartRem_5__3_), .B(
        n241), .CIN(rem_45_u_div_CryTmp_4__3_), .COUT(
        rem_45_u_div_CryTmp_4__4_), .SUM(rem_45_u_div_SumTmp_4__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_5_3 ( .A(rem_45_u_div_PartRem_6__3_), .B(
        n241), .CIN(rem_45_u_div_CryTmp_5__3_), .COUT(
        rem_45_u_div_CryTmp_5__4_), .SUM(rem_45_u_div_SumTmp_5__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_7_3 ( .A(rem_45_u_div_PartRem_8__3_), .B(
        n241), .CIN(rem_45_u_div_CryTmp_7__3_), .COUT(
        rem_45_u_div_CryTmp_7__4_), .SUM(rem_45_u_div_SumTmp_7__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_8_3 ( .A(rem_45_u_div_PartRem_9__3_), .B(
        n241), .CIN(rem_45_u_div_CryTmp_8__3_), .COUT(
        rem_45_u_div_CryTmp_8__4_), .SUM(rem_45_u_div_SumTmp_8__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_10_3 ( .A(rem_45_u_div_PartRem_11__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_10__3_), .COUT(
        rem_45_u_div_CryTmp_10__4_), .SUM(rem_45_u_div_SumTmp_10__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_11_3 ( .A(rem_45_u_div_PartRem_12__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_11__3_), .COUT(
        rem_45_u_div_CryTmp_11__4_), .SUM(rem_45_u_div_SumTmp_11__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_13_3 ( .A(rem_45_u_div_PartRem_14__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_13__3_), .COUT(
        rem_45_u_div_CryTmp_13__4_), .SUM(rem_45_u_div_SumTmp_13__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_14_3 ( .A(rem_45_u_div_PartRem_15__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_14__3_), .COUT(
        rem_45_u_div_CryTmp_14__4_), .SUM(rem_45_u_div_SumTmp_14__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_23_3 ( .A(rem_45_u_div_PartRem_24__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_23__3_), .COUT(
        rem_45_u_div_CryTmp_23__4_), .SUM(rem_45_u_div_SumTmp_23__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_6_3 ( .A(rem_45_u_div_PartRem_7__3_), .B(
        n241), .CIN(rem_45_u_div_CryTmp_6__3_), .COUT(
        rem_45_u_div_CryTmp_6__4_), .SUM(rem_45_u_div_SumTmp_6__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_9_3 ( .A(rem_45_u_div_PartRem_10__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_9__3_), .COUT(
        rem_45_u_div_CryTmp_9__4_), .SUM(rem_45_u_div_SumTmp_9__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_12_3 ( .A(rem_45_u_div_PartRem_13__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_12__3_), .COUT(
        rem_45_u_div_CryTmp_12__4_), .SUM(rem_45_u_div_SumTmp_12__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_15_3 ( .A(rem_45_u_div_PartRem_16__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_15__3_), .COUT(
        rem_45_u_div_CryTmp_15__4_), .SUM(rem_45_u_div_SumTmp_15__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_28_3 ( .A(rem_45_u_div_PartRem_29__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_28__3_), .COUT(
        rem_45_u_div_CryTmp_28__4_), .SUM(rem_45_u_div_SumTmp_28__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_13_1 ( .A(rem_45_u_div_PartRem_14__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_13__1_), .COUT(
        rem_45_u_div_CryTmp_13__2_), .SUM(rem_45_u_div_SumTmp_13__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_14_1 ( .A(rem_45_u_div_PartRem_15__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_14__1_), .COUT(
        rem_45_u_div_CryTmp_14__2_), .SUM(rem_45_u_div_SumTmp_14__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_15_1 ( .A(rem_45_u_div_PartRem_16__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_15__1_), .COUT(
        rem_45_u_div_CryTmp_15__2_), .SUM(rem_45_u_div_SumTmp_15__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_16_1 ( .A(rem_45_u_div_PartRem_17__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_16__1_), .COUT(
        rem_45_u_div_CryTmp_16__2_), .SUM(rem_45_u_div_SumTmp_16__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_17_1 ( .A(rem_45_u_div_PartRem_18__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_17__1_), .COUT(
        rem_45_u_div_CryTmp_17__2_), .SUM(rem_45_u_div_SumTmp_17__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_18_1 ( .A(rem_45_u_div_PartRem_19__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_18__1_), .COUT(
        rem_45_u_div_CryTmp_18__2_), .SUM(rem_45_u_div_SumTmp_18__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_26_1 ( .A(rem_45_u_div_PartRem_27__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_26__1_), .COUT(
        rem_45_u_div_CryTmp_26__2_), .SUM(rem_45_u_div_SumTmp_26__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_27_1 ( .A(rem_45_u_div_PartRem_28__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_27__1_), .COUT(
        rem_45_u_div_CryTmp_27__2_), .SUM(rem_45_u_div_SumTmp_27__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_28_1 ( .A(rem_45_u_div_PartRem_29__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_28__1_), .COUT(
        rem_45_u_div_CryTmp_28__2_), .SUM(rem_45_u_div_SumTmp_28__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_29_1 ( .A(rem_45_u_div_PartRem_30__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_29__1_), .COUT(
        rem_45_u_div_CryTmp_29__2_), .SUM(rem_45_u_div_SumTmp_29__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_13_2 ( .A(rem_45_u_div_PartRem_14__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_13__2_), .COUT(
        rem_45_u_div_CryTmp_13__3_), .SUM(rem_45_u_div_SumTmp_13__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_14_2 ( .A(rem_45_u_div_PartRem_15__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_14__2_), .COUT(
        rem_45_u_div_CryTmp_14__3_), .SUM(rem_45_u_div_SumTmp_14__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_15_2 ( .A(rem_45_u_div_PartRem_16__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_15__2_), .COUT(
        rem_45_u_div_CryTmp_15__3_), .SUM(rem_45_u_div_SumTmp_15__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_16_2 ( .A(rem_45_u_div_PartRem_17__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_16__2_), .COUT(
        rem_45_u_div_CryTmp_16__3_), .SUM(rem_45_u_div_SumTmp_16__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_17_2 ( .A(rem_45_u_div_PartRem_18__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_17__2_), .COUT(
        rem_45_u_div_CryTmp_17__3_), .SUM(rem_45_u_div_SumTmp_17__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_18_2 ( .A(rem_45_u_div_PartRem_19__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_18__2_), .COUT(
        rem_45_u_div_CryTmp_18__3_), .SUM(rem_45_u_div_SumTmp_18__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_27_2 ( .A(rem_45_u_div_PartRem_28__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_27__2_), .COUT(
        rem_45_u_div_CryTmp_27__3_), .SUM(rem_45_u_div_SumTmp_27__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_28_2 ( .A(rem_45_u_div_PartRem_29__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_28__2_), .COUT(
        rem_45_u_div_CryTmp_28__3_), .SUM(rem_45_u_div_SumTmp_28__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_1_3 ( .A(rem_45_u_div_PartRem_2__3_), .B(
        n241), .CIN(rem_45_u_div_CryTmp_1__3_), .COUT(
        rem_45_u_div_CryTmp_1__4_), .SUM(rem_45_u_div_SumTmp_1__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_19_2 ( .A(rem_45_u_div_PartRem_20__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_19__2_), .COUT(
        rem_45_u_div_CryTmp_19__3_), .SUM(rem_45_u_div_SumTmp_19__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_2_3 ( .A(rem_45_u_div_PartRem_3__3_), .B(
        n241), .CIN(rem_45_u_div_CryTmp_2__3_), .COUT(
        rem_45_u_div_CryTmp_2__4_), .SUM(rem_45_u_div_SumTmp_2__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_16_3 ( .A(rem_45_u_div_PartRem_17__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_16__3_), .COUT(
        rem_45_u_div_CryTmp_16__4_), .SUM(rem_45_u_div_SumTmp_16__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_17_3 ( .A(rem_45_u_div_PartRem_18__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_17__3_), .COUT(
        rem_45_u_div_CryTmp_17__4_), .SUM(rem_45_u_div_SumTmp_17__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_19_3 ( .A(rem_45_u_div_PartRem_20__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_19__3_), .COUT(
        rem_45_u_div_CryTmp_19__4_), .SUM(rem_45_u_div_SumTmp_19__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_22_1 ( .A(rem_45_u_div_PartRem_23__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_22__1_), .COUT(
        rem_45_u_div_CryTmp_22__2_), .SUM(rem_45_u_div_SumTmp_22__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_19_1 ( .A(rem_45_u_div_PartRem_20__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_19__1_), .COUT(
        rem_45_u_div_CryTmp_19__2_), .SUM(rem_45_u_div_SumTmp_19__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_20_1 ( .A(rem_45_u_div_PartRem_21__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_20__1_), .COUT(
        rem_45_u_div_CryTmp_20__2_), .SUM(rem_45_u_div_SumTmp_20__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_21_1 ( .A(rem_45_u_div_PartRem_22__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_21__1_), .COUT(
        rem_45_u_div_CryTmp_21__2_), .SUM(rem_45_u_div_SumTmp_21__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_23_1 ( .A(rem_45_u_div_PartRem_24__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_23__1_), .COUT(
        rem_45_u_div_CryTmp_23__2_), .SUM(rem_45_u_div_SumTmp_23__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_24_1 ( .A(rem_45_u_div_PartRem_25__1_), 
        .B(n243), .CIN(rem_45_u_div_CryTmp_24__1_), .COUT(
        rem_45_u_div_CryTmp_24__2_), .SUM(rem_45_u_div_SumTmp_24__1_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_20_2 ( .A(rem_45_u_div_PartRem_21__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_20__2_), .COUT(
        rem_45_u_div_CryTmp_20__3_), .SUM(rem_45_u_div_SumTmp_20__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_21_2 ( .A(rem_45_u_div_PartRem_22__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_21__2_), .COUT(
        rem_45_u_div_CryTmp_21__3_), .SUM(rem_45_u_div_SumTmp_21__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_22_2 ( .A(rem_45_u_div_PartRem_23__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_22__2_), .COUT(
        rem_45_u_div_CryTmp_22__3_), .SUM(rem_45_u_div_SumTmp_22__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_23_2 ( .A(rem_45_u_div_PartRem_24__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_23__2_), .COUT(
        rem_45_u_div_CryTmp_23__3_), .SUM(rem_45_u_div_SumTmp_23__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_24_2 ( .A(rem_45_u_div_PartRem_25__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_24__2_), .COUT(
        rem_45_u_div_CryTmp_24__3_), .SUM(rem_45_u_div_SumTmp_24__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_26_2 ( .A(rem_45_u_div_PartRem_27__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_26__2_), .COUT(
        rem_45_u_div_CryTmp_26__3_), .SUM(rem_45_u_div_SumTmp_26__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_20_3 ( .A(rem_45_u_div_PartRem_21__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_20__3_), .COUT(
        rem_45_u_div_CryTmp_20__4_), .SUM(rem_45_u_div_SumTmp_20__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_22_3 ( .A(rem_45_u_div_PartRem_23__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_22__3_), .COUT(
        rem_45_u_div_CryTmp_22__4_), .SUM(rem_45_u_div_SumTmp_22__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_25_3 ( .A(rem_45_u_div_PartRem_26__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_25__3_), .COUT(
        rem_45_u_div_CryTmp_25__4_), .SUM(rem_45_u_div_SumTmp_25__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_26_3 ( .A(rem_45_u_div_PartRem_27__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_26__3_), .COUT(
        rem_45_u_div_CryTmp_26__4_), .SUM(rem_45_u_div_SumTmp_26__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_29_2 ( .A(rem_45_u_div_PartRem_30__2_), 
        .B(n242), .CIN(rem_45_u_div_CryTmp_29__2_), .COUT(
        rem_45_u_div_CryTmp_29__3_), .SUM(rem_45_u_div_SumTmp_29__2_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_0_3 ( .A(rem_45_u_div_PartRem_1__3_), .B(
        n241), .CIN(rem_45_u_div_CryTmp_0__3_), .COUT(
        rem_45_u_div_CryTmp_0__4_), .SUM(rem_45_u_div_SumTmp_0__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_3_3 ( .A(rem_45_u_div_PartRem_4__3_), .B(
        n241), .CIN(rem_45_u_div_CryTmp_3__3_), .COUT(
        rem_45_u_div_CryTmp_3__4_), .SUM(rem_45_u_div_SumTmp_3__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_18_3 ( .A(rem_45_u_div_PartRem_19__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_18__3_), .COUT(
        rem_45_u_div_CryTmp_18__4_), .SUM(rem_45_u_div_SumTmp_18__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_21_3 ( .A(rem_45_u_div_PartRem_22__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_21__3_), .COUT(
        rem_45_u_div_CryTmp_21__4_), .SUM(rem_45_u_div_SumTmp_21__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_24_3 ( .A(rem_45_u_div_PartRem_25__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_24__3_), .COUT(
        rem_45_u_div_CryTmp_24__4_), .SUM(rem_45_u_div_SumTmp_24__3_) );
  ADDF_E rem_45_u_div_u_fa_PartRem_0_27_3 ( .A(rem_45_u_div_PartRem_28__3_), 
        .B(n241), .CIN(rem_45_u_div_CryTmp_27__3_), .COUT(
        rem_45_u_div_CryTmp_27__4_), .SUM(rem_45_u_div_SumTmp_27__3_) );
  DFF_E counter_reg_13_ ( .D(N71), .CLK(CLK_500K), .Q(n216), .QBAR(n434) );
  DFF_E counter_reg_12_ ( .D(N70), .CLK(CLK_500K), .Q(), .QBAR(n550) );
  DFF_E counter_reg_11_ ( .D(N69), .CLK(CLK_500K), .Q(n213), .QBAR(n540) );
  DFF_E counter_reg_10_ ( .D(N68), .CLK(CLK_500K), .Q(n211), .QBAR(n423) );
  DFF_E counter_reg_9_ ( .D(N67), .CLK(CLK_500K), .Q(n209), .QBAR(n53) );
  DFF_E counter_reg_8_ ( .D(N66), .CLK(CLK_500K), .Q(), .QBAR(n52) );
  DFF_E counter_reg_7_ ( .D(N65), .CLK(CLK_500K), .Q(n198), .QBAR(n51) );
  DFF_E counter_reg_6_ ( .D(N64), .CLK(CLK_500K), .Q(), .QBAR(n50) );
  DFF_E counter_reg_5_ ( .D(N63), .CLK(CLK_500K), .Q(n206), .QBAR(n49) );
  DFF_E counter_reg_4_ ( .D(N62), .CLK(CLK_500K), .Q(), .QBAR(n48) );
  DFF_E counter_reg_3_ ( .D(N61), .CLK(CLK_500K), .Q(n201), .QBAR(n47) );
  DFF_E counter_reg_1_ ( .D(N59), .CLK(CLK_500K), .Q(n205), .QBAR(n433) );
  DFF_E counter_reg_0_ ( .D(N58), .CLK(CLK_500K), .Q(n204), .QBAR(n440) );
  DFF_E counter_reg_14_ ( .D(N72), .CLK(CLK_500K), .Q(n218), .QBAR(n424) );
  DFF_E counter_reg_15_ ( .D(N73), .CLK(CLK_500K), .Q(n220), .QBAR(n56) );
  DFF_E counter_reg_2_ ( .D(N60), .CLK(CLK_500K), .Q(n202), .QBAR(n432) );
  DFF_E counter_reg_16_ ( .D(N74), .CLK(CLK_500K), .Q(n222), .QBAR(n57) );
  DFF_E counter_reg_18_ ( .D(N76), .CLK(CLK_500K), .Q(n226), .QBAR(n426) );
  DFF_E counter_reg_17_ ( .D(N75), .CLK(CLK_500K), .Q(n224), .QBAR(n425) );
  DFF_E VSTIM_P_Q_reg ( .D(N55), .CLK(CLK_500K), .Q(VSTIM_P), .QBAR() );
  DFF_E VSTIM_N_Q_reg ( .D(N54), .CLK(CLK_500K), .Q(VSTIM_N), .QBAR() );
  DFF_E DO_SAMPLE_Q_reg ( .D(n250), .CLK(CLK_500K), .Q(DO_SAMPLE), .QBAR(n170)
         );
  DFF_K MEASURE_PRESCALAR_Q_reg_3_ ( .D(MEASURE_PRESCALAR[3]), .CLK(CLK_500K), 
        .Q(), .QBAR(n241) );
  DFF_K MEASURE_PRESCALAR_Q_reg_2_ ( .D(MEASURE_PRESCALAR[2]), .CLK(CLK_500K), 
        .Q(), .QBAR(n242) );
  DFF_K MEASURE_PRESCALAR_Q_reg_1_ ( .D(MEASURE_PRESCALAR[1]), .CLK(CLK_500K), 
        .Q(), .QBAR(n243) );
  DFF_K MEASURE_PRESCALAR_Q_reg_0_ ( .D(MEASURE_PRESCALAR[0]), .CLK(CLK_500K), 
        .Q(n43), .QBAR(n441) );
  AO22_F U274 ( .A1(rem_45_u_div_SumTmp_30__1_), .A2(n240), .B1(1'b0), .B2(
        n354), .Z(rem_45_u_div_PartRem_30__2_) );
  INVERTBAL_H U420 ( .A(n43), .Z(rem_45_u_div_CryTmp_30__1_) );
  OAI21_C U421 ( .A1(rem_45_u_div_CryTmp_30__1_), .A2(n354), .B(1'b1), .Z(
        rem_45_u_div_PartRem_30__1_) );
  INVERTBAL_H U422 ( .A(n438), .Z(rem_45_u_div_CryTmp_29__1_) );
  OAI21_C U423 ( .A1(rem_45_u_div_CryTmp_29__1_), .A2(n351), .B(1'b1), .Z(
        rem_45_u_div_PartRem_29__1_) );
  INVERTBAL_H U424 ( .A(n438), .Z(rem_45_u_div_CryTmp_28__1_) );
  OAI21_C U425 ( .A1(rem_45_u_div_CryTmp_28__1_), .A2(n238), .B(1'b1), .Z(
        rem_45_u_div_PartRem_28__1_) );
  INVERTBAL_H U426 ( .A(n438), .Z(rem_45_u_div_CryTmp_27__1_) );
  OAI21_C U427 ( .A1(rem_45_u_div_CryTmp_27__1_), .A2(n237), .B(1'b1), .Z(
        rem_45_u_div_PartRem_27__1_) );
  INVERTBAL_H U428 ( .A(n437), .Z(rem_45_u_div_CryTmp_26__1_) );
  OAI21_C U429 ( .A1(rem_45_u_div_CryTmp_26__1_), .A2(n342), .B(1'b1), .Z(
        rem_45_u_div_PartRem_26__1_) );
  INVERTBAL_H U430 ( .A(n437), .Z(rem_45_u_div_CryTmp_25__1_) );
  OAI21_C U431 ( .A1(rem_45_u_div_CryTmp_25__1_), .A2(n338), .B(1'b1), .Z(
        rem_45_u_div_PartRem_25__1_) );
  INVERTBAL_H U432 ( .A(n437), .Z(rem_45_u_div_CryTmp_24__1_) );
  OAI21_C U433 ( .A1(rem_45_u_div_CryTmp_24__1_), .A2(n234), .B(1'b1), .Z(
        rem_45_u_div_PartRem_24__1_) );
  INVERTBAL_H U434 ( .A(n437), .Z(rem_45_u_div_CryTmp_23__1_) );
  OAI21_C U435 ( .A1(rem_45_u_div_CryTmp_23__1_), .A2(n331), .B(1'b1), .Z(
        rem_45_u_div_PartRem_23__1_) );
  INVERTBAL_H U436 ( .A(n437), .Z(rem_45_u_div_CryTmp_22__1_) );
  OAI21_C U437 ( .A1(rem_45_u_div_CryTmp_22__1_), .A2(n328), .B(1'b1), .Z(
        rem_45_u_div_PartRem_22__1_) );
  INVERTBAL_H U438 ( .A(n437), .Z(rem_45_u_div_CryTmp_21__1_) );
  OAI21_C U439 ( .A1(rem_45_u_div_CryTmp_21__1_), .A2(n231), .B(1'b1), .Z(
        rem_45_u_div_PartRem_21__1_) );
  INVERTBAL_H U440 ( .A(n437), .Z(rem_45_u_div_CryTmp_20__1_) );
  OAI21_C U441 ( .A1(rem_45_u_div_CryTmp_20__1_), .A2(n321), .B(1'b1), .Z(
        rem_45_u_div_PartRem_20__1_) );
  INVERTBAL_H U442 ( .A(n396), .Z(n361) );
  INVERTBAL_H U443 ( .A(n437), .Z(rem_45_u_div_CryTmp_19__1_) );
  OAI21_C U444 ( .A1(rem_45_u_div_CryTmp_19__1_), .A2(n318), .B(1'b1), .Z(
        rem_45_u_div_PartRem_19__1_) );
  OR4_E U445 ( .A(n414), .B(n211), .C(1'b0), .D(1'b0), .Z(n406) );
  AND2_F U446 ( .A(n243), .B(rem_45_u_div_CryTmp_30__1_), .Z(
        rem_45_u_div_CryTmp_30__2_) );
  XOR2_C U447 ( .A(rem_45_u_div_CryTmp_30__1_), .B(n243), .Z(
        rem_45_u_div_SumTmp_30__1_) );
  NOR4_B U448 ( .A(n422), .B(n220), .C(1'b0), .D(1'b0), .Z(n421) );
  AOI21_C U450 ( .A1(n223), .A2(rem_45_u_div_SumTmp_17__3_), .B(n320), .Z(n308) );
  AOI21_C U451 ( .A1(n317), .A2(rem_45_u_div_SumTmp_18__3_), .B(n323), .Z(n311) );
  AOI21_C U452 ( .A1(n229), .A2(rem_45_u_div_SumTmp_20__3_), .B(n330), .Z(n318) );
  AOI21_C U453 ( .A1(n192), .A2(rem_45_u_div_SumTmp_2__3_), .B(n267), .Z(n257)
         );
  AOI21_C U454 ( .A1(n264), .A2(rem_45_u_div_SumTmp_3__3_), .B(n271), .Z(n259)
         );
  AOI21_C U455 ( .A1(n236), .A2(rem_45_u_div_SumTmp_26__3_), .B(n350), .Z(n338) );
  AOI21_C U456 ( .A1(n325), .A2(rem_45_u_div_SumTmp_21__3_), .B(n333), .Z(n321) );
  NAND2_F U457 ( .A(n347), .B(n348), .Z(n335) );
  NAND2_F U458 ( .A(rem_45_u_div_SumTmp_25__3_), .B(n235), .Z(n348) );
  AOI21_C U459 ( .A1(n338), .A2(rem_45_u_div_PartRem_26__3_), .B(
        rem_45_u_div_CryTmp_24__4_), .Z(n347) );
  NAND2_F U460 ( .A(n336), .B(n337), .Z(n325) );
  NAND2_F U461 ( .A(rem_45_u_div_SumTmp_22__3_), .B(n232), .Z(n337) );
  AOI21_C U462 ( .A1(n328), .A2(rem_45_u_div_PartRem_23__3_), .B(
        rem_45_u_div_CryTmp_21__4_), .Z(n336) );
  NAND2_F U463 ( .A(n262), .B(n263), .Z(n256) );
  NAND2_F U464 ( .A(rem_45_u_div_SumTmp_1__3_), .B(n191), .Z(n263) );
  AOI21_C U465 ( .A1(n257), .A2(rem_45_u_div_PartRem_2__3_), .B(
        rem_45_u_div_CryTmp_0__4_), .Z(n262) );
  NAND2_F U466 ( .A(n326), .B(n327), .Z(n317) );
  NAND2_F U467 ( .A(rem_45_u_div_SumTmp_19__3_), .B(n227), .Z(n327) );
  AOI21_C U468 ( .A1(n318), .A2(rem_45_u_div_PartRem_20__3_), .B(
        rem_45_u_div_CryTmp_18__4_), .Z(n326) );
  AOI21_C U469 ( .A1(n346), .A2(rem_45_u_div_SumTmp_27__3_), .B(n353), .Z(n342) );
  AOI21_C U470 ( .A1(n217), .A2(rem_45_u_div_SumTmp_14__3_), .B(n310), .Z(n297) );
  AOI21_C U471 ( .A1(n212), .A2(rem_45_u_div_SumTmp_11__3_), .B(n299), .Z(n286) );
  AOI21_C U472 ( .A1(n207), .A2(rem_45_u_div_SumTmp_8__3_), .B(n288), .Z(n276)
         );
  AOI21_C U473 ( .A1(n273), .A2(rem_45_u_div_SumTmp_6__3_), .B(n281), .Z(n268)
         );
  AOI21_C U474 ( .A1(n294), .A2(rem_45_u_div_SumTmp_12__3_), .B(n303), .Z(n289) );
  AOI21_C U475 ( .A1(n307), .A2(rem_45_u_div_SumTmp_15__3_), .B(n313), .Z(n301) );
  AOI21_C U476 ( .A1(n233), .A2(rem_45_u_div_SumTmp_23__3_), .B(n341), .Z(n328) );
  AOI21_C U477 ( .A1(n195), .A2(rem_45_u_div_SumTmp_5__3_), .B(n278), .Z(n265)
         );
  AOI21_C U478 ( .A1(n285), .A2(rem_45_u_div_SumTmp_9__3_), .B(n292), .Z(n279)
         );
  NAND2_F U479 ( .A(n283), .B(n284), .Z(n273) );
  NAND2_F U480 ( .A(rem_45_u_div_SumTmp_7__3_), .B(n197), .Z(n284) );
  AOI21_C U481 ( .A1(n276), .A2(rem_45_u_div_PartRem_8__3_), .B(
        rem_45_u_div_CryTmp_6__4_), .Z(n283) );
  NAND2_F U482 ( .A(n305), .B(n306), .Z(n294) );
  NAND2_F U483 ( .A(rem_45_u_div_SumTmp_13__3_), .B(n215), .Z(n306) );
  AOI21_C U484 ( .A1(n297), .A2(rem_45_u_div_PartRem_14__3_), .B(
        rem_45_u_div_CryTmp_12__4_), .Z(n305) );
  NAND3_E U485 ( .A(n241), .B(n242), .C(rem_45_u_div_CryTmp_30__2_), .Z(n354)
         );
  OAI21_C U486 ( .A1(rem_45_u_div_CryTmp_1__1_), .A2(n257), .B(n258), .Z(
        rem_45_u_div_PartRem_1__1_) );
  OAI21_C U487 ( .A1(n257), .A2(n439), .B(n205), .Z(n258) );
  NAND2_F U488 ( .A(n295), .B(n296), .Z(n285) );
  NAND2_F U489 ( .A(rem_45_u_div_SumTmp_10__3_), .B(n210), .Z(n296) );
  AOI21_C U490 ( .A1(n286), .A2(rem_45_u_div_PartRem_11__3_), .B(
        rem_45_u_div_CryTmp_9__4_), .Z(n295) );
  NAND2_F U491 ( .A(n315), .B(n316), .Z(n307) );
  NAND2_F U492 ( .A(rem_45_u_div_SumTmp_16__3_), .B(n221), .Z(n316) );
  AOI21_C U493 ( .A1(n308), .A2(rem_45_u_div_PartRem_17__3_), .B(
        rem_45_u_div_CryTmp_15__4_), .Z(n315) );
  NAND2_F U494 ( .A(n274), .B(n275), .Z(n264) );
  NAND2_F U495 ( .A(rem_45_u_div_SumTmp_4__3_), .B(n194), .Z(n275) );
  AOI21_C U496 ( .A1(n265), .A2(rem_45_u_div_PartRem_5__3_), .B(
        rem_45_u_div_CryTmp_3__4_), .Z(n274) );
  NAND2_F U497 ( .A(rem_45_u_div_CryTmp_29__3_), .B(n241), .Z(n351) );
  OAI21_C U498 ( .A1(rem_45_u_div_CryTmp_10__1_), .A2(n286), .B(n287), .Z(
        rem_45_u_div_PartRem_10__1_) );
  OAI21_C U499 ( .A1(n286), .A2(n441), .B(n211), .Z(n287) );
  OAI21_C U500 ( .A1(rem_45_u_div_CryTmp_11__1_), .A2(n289), .B(n291), .Z(
        rem_45_u_div_PartRem_11__1_) );
  OAI21_C U501 ( .A1(n289), .A2(n439), .B(n213), .Z(n291) );
  OAI21_C U502 ( .A1(rem_45_u_div_CryTmp_5__1_), .A2(n268), .B(n269), .Z(
        rem_45_u_div_PartRem_5__1_) );
  OAI21_C U503 ( .A1(n268), .A2(n439), .B(n206), .Z(n269) );
  OAI21_C U504 ( .A1(rem_45_u_div_CryTmp_2__1_), .A2(n259), .B(n260), .Z(
        rem_45_u_div_PartRem_2__1_) );
  OAI21_C U505 ( .A1(n259), .A2(n441), .B(n202), .Z(n260) );
  OAI21_C U506 ( .A1(rem_45_u_div_CryTmp_18__1_), .A2(n225), .B(n314), .Z(
        rem_45_u_div_PartRem_18__1_) );
  OAI21_C U507 ( .A1(n225), .A2(n439), .B(n226), .Z(n314) );
  OAI21_C U508 ( .A1(rem_45_u_div_CryTmp_9__1_), .A2(n208), .B(n282), .Z(
        rem_45_u_div_PartRem_9__1_) );
  OAI21_C U509 ( .A1(n208), .A2(n441), .B(n209), .Z(n282) );
  OAI21_C U510 ( .A1(rem_45_u_div_CryTmp_3__1_), .A2(n193), .B(n261), .Z(
        rem_45_u_div_PartRem_3__1_) );
  OAI21_C U511 ( .A1(n193), .A2(n441), .B(n201), .Z(n261) );
  OAI21_C U512 ( .A1(rem_45_u_div_CryTmp_15__1_), .A2(n219), .B(n304), .Z(
        rem_45_u_div_PartRem_15__1_) );
  OAI21_C U513 ( .A1(n219), .A2(n439), .B(n220), .Z(n304) );
  NAND2_F U514 ( .A(n356), .B(n357), .Z(n346) );
  NAND2_F U515 ( .A(rem_45_u_div_SumTmp_28__3_), .B(rem_45_u_div_CryTmp_28__4_), .Z(n357) );
  AOI21_C U516 ( .A1(rem_45_u_div_PartRem_29__3_), .A2(n238), .B(
        rem_45_u_div_CryTmp_27__4_), .Z(n356) );
  OAI21_C U517 ( .A1(rem_45_u_div_CryTmp_7__1_), .A2(n276), .B(n277), .Z(
        rem_45_u_div_PartRem_7__1_) );
  OAI21_C U518 ( .A1(n276), .A2(n439), .B(n198), .Z(n277) );
  OAI21_C U519 ( .A1(rem_45_u_div_CryTmp_13__1_), .A2(n297), .B(n298), .Z(
        rem_45_u_div_PartRem_13__1_) );
  OAI21_C U520 ( .A1(n297), .A2(n439), .B(n216), .Z(n298) );
  OAI21_C U521 ( .A1(rem_45_u_div_CryTmp_16__1_), .A2(n308), .B(n309), .Z(
        rem_45_u_div_PartRem_16__1_) );
  OAI21_C U522 ( .A1(n308), .A2(n439), .B(n222), .Z(n309) );
  OAI21_C U523 ( .A1(rem_45_u_div_CryTmp_14__1_), .A2(n301), .B(n302), .Z(
        rem_45_u_div_PartRem_14__1_) );
  OAI21_C U524 ( .A1(n301), .A2(n439), .B(n218), .Z(n302) );
  OAI21_C U525 ( .A1(rem_45_u_div_CryTmp_17__1_), .A2(n311), .B(n312), .Z(
        rem_45_u_div_PartRem_17__1_) );
  OAI21_C U526 ( .A1(n311), .A2(n439), .B(n224), .Z(n312) );
  AOI21_C U527 ( .A1(n335), .A2(rem_45_u_div_SumTmp_24__3_), .B(n344), .Z(n331) );
  OAI22_B U528 ( .A1(n190), .A2(n254), .B1(n255), .B2(n256), .Z(n253) );
  NOR4_B U529 ( .A(rem_45_u_div_PartRem_1__3_), .B(rem_45_u_div_PartRem_1__2_), 
        .C(rem_45_u_div_PartRem_1__1_), .D(n204), .Z(n255) );
  NOR4_B U530 ( .A(rem_45_u_div_SumTmp_0__3_), .B(rem_45_u_div_SumTmp_0__2_), 
        .C(rem_45_u_div_SumTmp_0__1_), .D(n247), .Z(n254) );
  INVERT_I U531 ( .A(n441), .Z(n438) );
  INVERT_I U532 ( .A(n439), .Z(n437) );
  NAND2_F U533 ( .A(n378), .B(n209), .Z(n376) );
  NAND2_F U534 ( .A(n391), .B(n201), .Z(n389) );
  NAND2_F U535 ( .A(n374), .B(n213), .Z(n372) );
  NAND2_F U536 ( .A(n387), .B(n206), .Z(n385) );
  NAND2_F U537 ( .A(n370), .B(n216), .Z(n368) );
  NAND2_F U538 ( .A(n366), .B(n220), .Z(n364) );
  NAND2_F U539 ( .A(n383), .B(n198), .Z(n381) );
  NOR2_E U540 ( .A(n436), .B(n363), .Z(N75) );
  NOR2_E U541 ( .A(n436), .B(n367), .Z(N73) );
  NOR2_E U542 ( .A(n436), .B(n371), .Z(N71) );
  NAND2_F U543 ( .A(n416), .B(n206), .Z(n408) );
  NOR2_E U544 ( .A(n436), .B(n204), .Z(N58) );
  NOR2_E U545 ( .A(n436), .B(n379), .Z(N67) );
  NOR2_E U546 ( .A(n436), .B(n392), .Z(N61) );
  NOR2_E U547 ( .A(n436), .B(n375), .Z(N69) );
  NOR2_E U548 ( .A(n395), .B(n436), .Z(N59) );
  NOR2_E U549 ( .A(n436), .B(n388), .Z(N63) );
  NOR2_E U550 ( .A(n436), .B(n384), .Z(N65) );
  OAI21_C U551 ( .A1(rem_45_u_div_CryTmp_4__1_), .A2(n265), .B(n266), .Z(
        rem_45_u_div_PartRem_4__1_) );
  OAI21_C U552 ( .A1(rem_45_u_div_CryTmp_12__1_), .A2(n214), .B(n293), .Z(
        rem_45_u_div_PartRem_12__1_) );
  OAI21_C U553 ( .A1(rem_45_u_div_CryTmp_6__1_), .A2(n196), .B(n272), .Z(
        rem_45_u_div_PartRem_6__1_) );
  OAI21_C U554 ( .A1(rem_45_u_div_CryTmp_8__1_), .A2(n279), .B(n280), .Z(
        rem_45_u_div_PartRem_8__1_) );
  OAI22_B U555 ( .A1(n170), .A2(n248), .B1(DO_SAMPLE), .B2(n249), .Z(n250) );
  NAND2_F U556 ( .A(n248), .B(n251), .Z(n249) );
  OAI21_C U557 ( .A1(n252), .A2(n253), .B(n251), .Z(n248) );
  INVERT_I U558 ( .A(n43), .Z(n439) );
  NAND2_F U559 ( .A(n426), .B(n437), .Z(rem_45_u_div_CryTmp_18__1_) );
  NAND2_F U560 ( .A(n425), .B(n437), .Z(rem_45_u_div_CryTmp_17__1_) );
  NAND2_F U561 ( .A(n57), .B(n437), .Z(rem_45_u_div_CryTmp_16__1_) );
  NAND2_F U562 ( .A(n56), .B(n437), .Z(rem_45_u_div_CryTmp_15__1_) );
  NAND2_F U563 ( .A(n424), .B(n437), .Z(rem_45_u_div_CryTmp_14__1_) );
  NAND2_F U564 ( .A(n434), .B(n43), .Z(rem_45_u_div_CryTmp_13__1_) );
  NAND2_F U565 ( .A(n550), .B(n43), .Z(rem_45_u_div_CryTmp_12__1_) );
  NAND2_F U566 ( .A(n540), .B(n43), .Z(rem_45_u_div_CryTmp_11__1_) );
  NAND2_F U567 ( .A(n423), .B(n43), .Z(rem_45_u_div_CryTmp_10__1_) );
  NAND2_F U568 ( .A(n53), .B(n43), .Z(rem_45_u_div_CryTmp_9__1_) );
  NAND2_F U569 ( .A(n52), .B(n43), .Z(rem_45_u_div_CryTmp_8__1_) );
  NAND2_F U570 ( .A(n51), .B(n43), .Z(rem_45_u_div_CryTmp_7__1_) );
  NAND2_F U571 ( .A(n50), .B(n43), .Z(rem_45_u_div_CryTmp_6__1_) );
  NAND2_F U572 ( .A(n49), .B(n43), .Z(rem_45_u_div_CryTmp_5__1_) );
  NAND2_F U573 ( .A(n48), .B(n43), .Z(rem_45_u_div_CryTmp_4__1_) );
  NAND2_F U574 ( .A(n47), .B(n43), .Z(rem_45_u_div_CryTmp_3__1_) );
  NAND2_F U575 ( .A(n432), .B(n43), .Z(rem_45_u_div_CryTmp_2__1_) );
  NAND2_F U576 ( .A(n433), .B(n437), .Z(rem_45_u_div_CryTmp_1__1_) );
  NOR3_B U577 ( .A(n433), .B(n432), .C(n440), .Z(n391) );
  NOR2_E U578 ( .A(n389), .B(n48), .Z(n387) );
  NOR2_E U579 ( .A(n372), .B(n550), .Z(n370) );
  NOR2_E U580 ( .A(n385), .B(n50), .Z(n383) );
  NOR2_E U581 ( .A(n376), .B(n423), .Z(n374) );
  NOR2_E U582 ( .A(n381), .B(n52), .Z(n378) );
  NOR2_E U583 ( .A(n368), .B(n424), .Z(n366) );
  NOR2_E U584 ( .A(n364), .B(n57), .Z(n362) );
  NOR2_E U585 ( .A(n436), .B(n365), .Z(N74) );
  AOI21_C U586 ( .A1(n426), .A2(n359), .B(n436), .Z(N76) );
  NAND2_F U587 ( .A(n362), .B(n224), .Z(n359) );
  NOR2_E U588 ( .A(n204), .B(n439), .Z(n247) );
  NOR3_B U589 ( .A(n51), .B(n52), .C(n50), .Z(n416) );
  OAI21_C U590 ( .A1(n432), .A2(n393), .B(n394), .Z(N60) );
  NAND4_B U591 ( .A(n199), .B(n432), .C(n204), .D(n205), .Z(n394) );
  AOI21_C U592 ( .A1(n199), .A2(n433), .B(N58), .Z(n393) );
  BUFFER_I U593 ( .A(n361), .Z(n436) );
  OAI21_C U594 ( .A1(n222), .A2(n402), .B(n226), .Z(n396) );
  OAI21_C U595 ( .A1(n403), .A2(n56), .B(n425), .Z(n402) );
  NOR3_B U596 ( .A(n216), .B(n404), .C(n218), .Z(n403) );
  AOI21_C U597 ( .A1(n405), .A2(n423), .B(n550), .Z(n404) );
  AOI21_C U598 ( .A1(n200), .A2(n209), .B(n213), .Z(n405) );
  NOR2_E U599 ( .A(n436), .B(n369), .Z(N72) );
  NOR2_E U600 ( .A(n436), .B(n373), .Z(N70) );
  NOR2_E U601 ( .A(n436), .B(n390), .Z(N62) );
  NOR2_E U602 ( .A(n436), .B(n386), .Z(N64) );
  NOR2_E U603 ( .A(n436), .B(n382), .Z(N66) );
  NOR2_E U604 ( .A(n436), .B(n377), .Z(N68) );
  NAND3_E U605 ( .A(n415), .B(n408), .C(n53), .Z(n413) );
  NAND4_B U606 ( .A(n416), .B(n410), .C(n417), .D(n201), .Z(n415) );
  NAND4_B U607 ( .A(n550), .B(n434), .C(n420), .D(n421), .Z(n414) );
  NOR3_B U608 ( .A(n218), .B(n222), .C(n213), .Z(n420) );
  NAND2_F U609 ( .A(n425), .B(n426), .Z(n422) );
  NAND2_F U610 ( .A(n440), .B(n433), .Z(n410) );
  NOR2_E U611 ( .A(n432), .B(n48), .Z(n417) );
  NOR2_E U612 ( .A(n411), .B(n251), .Z(N54) );
  AOI21_C U613 ( .A1(n418), .A2(n200), .B(n406), .Z(n411) );
  AOI21_C U614 ( .A1(n47), .A2(n48), .B(n53), .Z(n418) );
  NOR2_E U615 ( .A(n440), .B(n43), .Z(n252) );
  NOR3_B U616 ( .A(n406), .B(n407), .C(n209), .Z(N55) );
  NOR3_B U617 ( .A(n408), .B(n48), .C(n409), .Z(n407) );
  AOI21_C U618 ( .A1(n410), .A2(n202), .B(n201), .Z(n409) );
endmodule
